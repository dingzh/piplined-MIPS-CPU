`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:38:14 02/27/2016 
// Design Name: 
// Module Name:    Top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Top(
    input CLOCK,
    input wire RESET,
	 input [2:0] MODE,
	 output [7:0] LED,
	 input FAST
    );
////          GENRERATING SLOW CLOCK            /////////////
	wire CLOCK_IN;
	reg [26:0] Buffer = 0;
	always@ (posedge CLOCK) Buffer = Buffer + 1;
	assign CLOCK_IN = FAST ? Buffer[1] : Buffer[0];

////				IO MODE SEL							//////////////
	assign LED[7] = RESET;
	assign LED[6] = CLOCK_IN;
	wire [5:0] OUTPUT;
	assign LED[5:0] = OUTPUT;
	wire [31:0] reg1;
	wire [31:0] reg2;
	wire [7:0]  reg12;
	assign reg12[5:3] = reg2;
	assign reg12[2:0] = reg1;
	wire [31:0] CURR_PC_IO;
	wire [5:0] TEMP1;
	wire [5:0] TEMP2;
	assign TEMP1 = MODE[0] ? reg1:reg12;
	assign TEMP2 = MODE[1] ? reg2:TEMP1;
	assign OUTPUT = MODE[2]? CURR_PC_IO>>2:TEMP2;


//////             main control signal              / /////
	wire REG_DST,
		  JUMP,
		  BRANCH,
		  MEM_READ,
		  MEM_TO_REG,
		  MEM_WRITE,
		  ALU_SRC,
		  REG_WRITE,
		  ZERO;  //generated by ALU
	wire [1:0]  ALU_OP;
	wire [3:0]  ALU_CTR;
	
/////////         data bus                        //////

	wire [31:0] REG_DATA_1;
	wire [31:0] REG_DATA_2;  //reg read output
	wire [4:0]  REG_WRITE_ADDRESS;//reg write address, the data will be from the MEM_REG_MUX
	wire [31:0] ALU_RES;
	wire [31:0] EXTENDED_RES;
	
	wire [31:0] MEM_READ_DATA;	//address specified by alu result
	
	wire [31:0] MEM_REG_MUX;	//to be written into reg(memomy or alu result)
	wire [31:0] REG_ALU_MUX;  //which one to be used by ALU as the 2nd src(rt or imm)
	
/////////////////////////////////////////////////////////////////////////////////////////
//Instruction Memory
/////////////////	////////////////////////////////////////////////////////////////////////
	reg [31:0] InstrMemory[9:0]; 
	initial $readmemb("./src/inst.txt",InstrMemory);
	//define AND initial Instruction Memory
	wire [31:0] INSTR;	
	wire [31:0] PCp4;
   wire [31:0] CURR_PC;
	assign CURR_PC_IO = CURR_PC; //for the output part
	assign INSTR = InstrMemory[CURR_PC>>2];  //fetch instruction by PC
	
/////////////////////////////////////////////////////////////////////////////////////////
//generating PC
/////////////////////////////////////////////////////////////////////////////////////////
	wire [31:0] JUMP_ADDRESS;
	wire [31:0] BEQ_ADDRESS;
	//assign JUMP_ADDRESS
	assign JUMP_ADDRESS[31:28] = PCp4[31:28];
	assign JUMP_ADDRESS[27:2]  = INSTR[25:0];
	assign JUMP_ADDRESS[1:0]   = 'b00;
	//assign BEQ_ADDRESS
	assign BEQ_ADDRESS[31:0] = (EXTENDED_RES<<2) + PCp4;	
	
	wire [31:0] PC_SRC_SEL;
   wire [31:0] NEXT_PC;
	//wire [31:0] PCp4;
	//wire [31:0] CURR_PC;  //declared above;
	wire PC_SRC;
	assign PC_SRC = BRANCH & ZERO;	
	assign PCp4[31:0] = CURR_PC[31:0] + 4;
	//serval MUX below
	assign PC_SRC_SEL[31:0] = PC_SRC ? BEQ_ADDRESS[31:0]: PCp4[31:0];
	assign NEXT_PC[31:0] = JUMP ? JUMP_ADDRESS[31:0] : PC_SRC_SEL[31:0];
	
	
	//serval MUX below:
	assign MEM_REG_MUX = MEM_TO_REG ? MEM_READ_DATA : ALU_RES;	//REG_WRITE_DATA
	//R-type or load word
	assign REG_ALU_MUX = ALU_SRC ? EXTENDED_RES : REG_DATA_2;  
	//which one to be used by ALU as the 2nd src
	assign REG_WRITE_ADDRESS = REG_DST ? INSTR[15:11] : INSTR[20:16];
	//which reg will be written
	
////////////////////////////////////////////////////////////////////////
//instances
////////////////////////////////////////////////////////////////////////	
	Pc mainPC(
      .clock_in(CLOCK_IN),
      .nextPC(NEXT_PC),
      .currPC(CURR_PC),
		.rst(RESET)
    );	
	
	Ctr mainCtr(
		.opCode(INSTR[31:26]), 
		.regDst(REG_DST), 
		.aluSrc(ALU_SRC), 
		.memToReg(MEM_TO_REG), 
		.regWrite(REG_WRITE), 
		.memRead(MEM_READ), 
		.memWrite(MEM_WRITE), 
		.branch(BRANCH), 
		.aluOp(ALU_OP), 
		.jump(JUMP)
	);
	
	AluCtr mainAluCtr (
		.aluOp(ALU_OP), 
		.funct(INSTR[5:0]), 
		.aluCtr(ALU_CTR)
	);
	
	Alu mainAlu (
		.input1(REG_DATA_1), 
		.input2(REG_ALU_MUX), 
		.aluCtr(ALU_CTR), 
		.zero(ZERO), 
		.aluRes(ALU_RES)
	);
	
	signExt mainSignExt (
		.inst(INSTR[15:0]),
		.data(EXTENDED_RES)
	);
	
	dataMemory mainDataMemory (
		.clock_in(CLOCK_IN), 
		.address(ALU_RES), 
		.writeData(REG_DATA_2), 
		.readData(MEM_READ_DATA), 
		.memWrite(MEM_WRITE), 
		.memRead(MEM_READ)
	);
	
	Register mainRegister (
		.clock_in(CLOCK_IN), 
		.regWrite(REG_WRITE), 
		.readReg1(INSTR[25:21]), 
		.readReg2(INSTR[20:16]), 
		.writeReg(REG_WRITE_ADDRESS), 
		.writeData(MEM_REG_MUX), 
		.reset(RESET),
		.readData1(REG_DATA_1), 
		.readData2(REG_DATA_2),
		.reg1(reg1),
		.reg2(reg2)
	);	
	
endmodule
